// Code your testbench here
// or browse Examples
module tb();
  
  
endmodule